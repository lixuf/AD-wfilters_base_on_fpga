module xiaobo_top(
);
endmodule

