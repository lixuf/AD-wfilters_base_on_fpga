module xiaobo_top(
output fifo_xb_rreq,
input [15:0] fifo_xb_r_data,
input [2:0]fifo_xb_use,//滞后一个时钟
input fifo_xb_full
);
endmodule
